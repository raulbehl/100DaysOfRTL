// Simple interface for a mux

interface day14_if ();

  logic [3:0] req;
  logic [3:0] gnt;

endinterface
