`include "riscv_fetch.sv"
`include "riscv_decode.sv"
`include "riscv_regfile.sv"
`include "riscv_execute.sv"

module riscv_top (
  input		wire		clk,
  input		wire		reset
);
  
  // Instantiate and connect all the submodules
  
endmodule
