// Simple interface for a mux

interface day4_if ();

  logic [7:0]   a;
  logic [7:0]   b;
  logic [2:0]   op;
  logic [7:0]   alu;

endinterface
