// Simple interface for a mux

interface day1_if ();

  logic [7:0] a;
  logic [7:0] b;
  logic       sel;
  logic [7:0] y;

endinterface
