// Hello world from SV classes

class day22;

  function new();
    // Nothing to do here
  endfunction

  function void print_hello();
    $display("Hello, World!\n");
  endfunction

endclass
