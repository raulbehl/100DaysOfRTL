interface riscv_reg_intf ();
  
  logic [31:0] regfile[31:0];
  
endinterface