// Code your testbench here
// or browse Examples
