`include "riscv_fetch.sv"
`include "riscv_decode.sv"

module riscv_top (
  input		wire		clk,
  input		wire		reset
);
  
  // Instantiate and connect all the submodules
  
endmodule